typedef 6  NumInputs;
typedef 20 CyclesResolution;
typedef 4  TimeStampBytes;

typedef 8 NumLeds;
typedef 1 Log2LedPersistence;
typedef 1 Log2ErrorBlink;

typedef 15 AddrSize;

Bit#(8) dacCalibCycles = 50;
