typedef 6  NumInputs;
typedef 50 CyclesResolution;
typedef 4  TimeStampBytes;

typedef 8  NumLeds;
typedef 13 Log2LedPersistence;
typedef 7  Log2ErrorBlink;

typedef 15 AddrSize;

Bit#(19) dacCalibCycles = 500000;  // 10 ms
